module primer

fn main() {
	println('Simple ECS implementation in V')
}
